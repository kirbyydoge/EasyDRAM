`define DQ_WIDTH 64
`define ODT_WIDTH 1
`define CS_WIDTH 1
`define CKE_WIDTH 1
`define CK_WIDTH 1
`define ROW_ADDR_WIDTH 17

